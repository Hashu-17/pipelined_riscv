
module top(input clk, input reset);
    // Instantiate all pipeline stages and connect them here
    // This file is meant to orchestrate the complete datapath and control path
endmodule
